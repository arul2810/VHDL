module clock(

input clock1,

input clock2,

input a,

output q

);


always @ (posedge clock1 ) begin


end

endmodule
